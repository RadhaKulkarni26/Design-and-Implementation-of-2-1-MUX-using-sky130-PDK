* c:\spb_data\esim-workspace\multiplexer\multiplexer.cir

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

xM1  Net-_M1-Pad1_ select vdd vdd sky130_fd_pr__pfet_01v8		
xM7  Net-_M1-Pad1_ select GND GND sky130_fd_pr__nfet_01v8		
xM6  vout Net-_M12-Pad2_ vdd vdd sky130_fd_pr__pfet_01v8		
xM12  vout Net-_M12-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
xM2  Net-_M2-Pad1_ vin_1 vdd vdd sky130_fd_pr__pfet_01v8		
xM4  Net-_M12-Pad2_ vin_2 Net-_M2-Pad1_ vdd sky130_fd_pr__pfet_01v8		
xM3  Net-_M2-Pad1_ Net-_M1-Pad1_ vdd vdd sky130_fd_pr__pfet_01v8		
xM5  Net-_M12-Pad2_ select Net-_M2-Pad1_ vdd sky130_fd_pr__pfet_01v8		
xM8  Net-_M12-Pad2_ vin_1 Net-_M10-Pad1_ GND sky130_fd_pr__nfet_01v8		
xM10  Net-_M10-Pad1_ Net-_M1-Pad1_ GND GND sky130_fd_pr__nfet_01v8		
xM9  Net-_M12-Pad2_ vin_2 Net-_M11-Pad1_ GND sky130_fd_pr__nfet_01v8		
xM11  Net-_M11-Pad1_ select GND GND sky130_fd_pr__nfet_01v8	

Vdd vdd 0 3	
Vin_1 vin_1 0 pulse(0 3 0s 0s 0s 5us 10us)
Vin_2 vin_2 0 pulse(0 3 0s 0s 0s 2.5us 5us) 
Vd0 select 0 pulse(3 0 0s 0s 0s 10us 20us) 

.tran 0.1us 40us
.control
run
plot V(vin_1) V(vin_2) V(select) V(vout)
.endc

.end	
